module ins_rom(addr,Data);
input[10:0] addr;
output[11:0] Data;
reg[11:0] Data;

always @(addr)
begin

case(addr)

'd00000: Data = 12'b101000000001;
'd00001: Data = 12'b000001100011;
'd00002: Data = 12'b000001100101;
'd00003: Data = 12'b000001100110;
'd00004: Data = 12'b110011111000;
'd00005: Data = 12'b000000000101;
'd00006: Data = 12'b110000000000;
'd00007: Data = 12'b000000000110;
'd00008: Data = 12'b000001100101;
'd00009: Data = 12'b100101001110;
'd00010: Data = 12'b110000111000;
'd00011: Data = 12'b100101000000;
'd00012: Data = 12'b110000000000;
'd00013: Data = 12'b111000000111;
'd00014: Data = 12'b110100001000;
'd00015: Data = 12'b100101000000;
'd00016: Data = 12'b110000000001;
'd00017: Data = 12'b100101000000;
'd00018: Data = 12'b110000000100;
'd00019: Data = 12'b111000000111;
'd00020: Data = 12'b110100001000;
'd00021: Data = 12'b100101000000;
'd00022: Data = 12'b110000000010;
'd00023: Data = 12'b111000000011;
'd00024: Data = 12'b110100000100;
'd00025: Data = 12'b100101000000;
'd00026: Data = 12'b110000110000;
'd00027: Data = 12'b000000110010;
'd00028: Data = 12'b110000000000;
'd00029: Data = 12'b110110000000;
'd00030: Data = 12'b100101000000;
'd00031: Data = 12'b110000000000;
'd00032: Data = 12'b000000110001;
'd00033: Data = 12'b100101010100;
'd00034: Data = 12'b111011111111;
'd00035: Data = 12'b011001000011;
'd00036: Data = 12'b101000101000;
'd00037: Data = 12'b100100110111;
'd00038: Data = 12'b001010010001;
'd00039: Data = 12'b101000100000;
'd00040: Data = 12'b101000101000;
'd00041: Data = 12'b110011111111;
'd00042: Data = 12'b000000000110;
'd00043: Data = 12'b010000000101;
'd00044: Data = 12'b010100100101;
'd00045: Data = 12'b010101000101;
'd00046: Data = 12'b001000000110;
'd00047: Data = 12'b010001000101;
'd00048: Data = 12'b111010000000;
'd00049: Data = 12'b011101000011;
'd00050: Data = 12'b101000101001;
'd00051: Data = 12'b010000100101;
'd00052: Data = 12'b110000000000;
'd00053: Data = 12'b000000000110;
'd00054: Data = 12'b100000000000;
'd00055: Data = 12'b000000110000;
'd00056: Data = 12'b100100101001;
'd00057: Data = 12'b010000100101;
'd00058: Data = 12'b010100000101;
'd00059: Data = 12'b010101000101;
'd00060: Data = 12'b001000010000;
'd00061: Data = 12'b000000100110;
'd00062: Data = 12'b010001000101;
'd00063: Data = 12'b100000000000;
'd00064: Data = 12'b000000110000;
'd00065: Data = 12'b100100101001;
'd00066: Data = 12'b010000100101;
'd00067: Data = 12'b010000000101;
'd00068: Data = 12'b010101000101;
'd00069: Data = 12'b001000010000;
'd00070: Data = 12'b000000100110;
'd00071: Data = 12'b010001000101;
'd00072: Data = 12'b100000000000;
'd00073: Data = 12'b110000000001;
'd00074: Data = 12'b000000110011;
'd00075: Data = 12'b001011110011;
'd00076: Data = 12'b101001001011;
'd00077: Data = 12'b100000000000;
'd00078: Data = 12'b110000000001;
'd00079: Data = 12'b000000110100;
'd00080: Data = 12'b100101001001;
'd00081: Data = 12'b001011110100;
'd00082: Data = 12'b101001010000;
'd00083: Data = 12'b100000000000;
'd00084: Data = 12'b000111100010;
'd00085: Data = 12'b100001001000;
'd00086: Data = 12'b100001100101;
'd00087: Data = 12'b100001101100;
'd00088: Data = 12'b100001101100;
'd00089: Data = 12'b100001101111;
'd00090: Data = 12'b100000100000;
'd00091: Data = 12'b100000000000;
 
default: Data = 12'b000000000000;

endcase
end

endmodule
